-- Add some new file, to see what happen in git