-- Try to git clone and push to a repo on github. 
-- Add some text